library IEEE;
use IEEE.std_logic_1164.all;

entity com3 is
end entity com3;

architecture RTL of com3 is
begin
end architecture RTL;
