library IEEE;
use IEEE.std_logic_1164.all;

package pkg2 is

   component com1 is
   --
   end component com1;

   component com3 is
   --
   end component com3;

end package pkg2;
