library IEEE;
use IEEE.std_logic_1164.all;

package pkg1 is

   component com1 is
   --
   end component com1;

   component com2 is
   --
   end component com2;

end package pkg1;
