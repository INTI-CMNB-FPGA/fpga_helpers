library IEEE;
use IEEE.std_logic_1164.all;

entity com5 is
end entity com5;

architecture RTL of com5 is
begin
end architecture RTL;
