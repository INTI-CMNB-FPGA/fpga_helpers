library IEEE;
use IEEE.std_logic_1164.all;

package pkg3 is

   component com5 is
   --
   end component com5;

end package pkg3;
