library IEEE;
use IEEE.std_logic_1164.all;

entity com2 is
end entity com2;

architecture RTL of com2 is
begin
end architecture RTL;
