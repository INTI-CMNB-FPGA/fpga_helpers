library IEEE;
use IEEE.std_logic_1164.all;

entity com4 is
end entity com4;

architecture RTL of com4 is
begin
end architecture RTL;
