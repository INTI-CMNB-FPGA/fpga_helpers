library IEEE;
use IEEE.std_logic_1164.all;

entity com1 is
end entity com1;

architecture RTL of com1 is
begin
end architecture RTL;
